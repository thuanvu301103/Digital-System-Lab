CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
280 130 6 290 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
176 438 1534 795
9437202 0
0
6 Title:
5 Name:
0
0
0
10
5 4081~
219 655 301 0 3 22
0 5 6 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
4983 0 0
2
44767.9 0
0
5 4071~
219 687 268 0 3 22
0 2 4 3
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3628 0 0
2
44767.9 0
0
2 +V
167 375 229 0 1 3
0 7
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4875 0 0
2
44767.9 0
0
14 Logic Display~
6 575 155 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8832 0 0
2
44767.9 0
0
14 Logic Display~
6 551 156 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3372 0 0
2
44767.9 0
0
14 Logic Display~
6 527 157 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
876 0 0
2
44767.9 0
0
14 Logic Display~
6 502 157 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 D
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5386 0 0
2
44767.9 0
0
7 Pulser~
4 311 286 0 10 12
0 13 14 12 15 0 0 10 10 10
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
890 0 0
2
44767.9 0
0
6 74LS73
102 571 285 0 12 25
0 7 7 9 3 7 7 10 3 10
5 11 2
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 0 0 0 0 0
1 U
3580 0 0
2
44767.9 0
0
6 74LS73
102 448 286 0 12 25
0 7 7 12 3 7 7 8 3 8
16 9 6
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 0 0 0 0
1 U
7445 0 0
2
44767.9 0
0
24
12 1 2 0 0 8320 0 9 2 0 0 3
609 312
609 259
674 259
8 0 3 0 0 4096 0 9 0 0 5 2
533 321
533 363
8 0 3 0 0 0 0 10 0 0 5 2
410 322
410 363
4 0 3 0 0 8192 0 9 0 0 5 3
533 285
512 285
512 363
3 4 3 0 0 8320 0 2 10 0 0 5
720 268
720 363
389 363
389 286
410 286
3 2 4 0 0 8320 0 1 2 0 0 4
676 301
675 301
675 277
674 277
10 1 5 0 0 4224 0 9 1 0 0 4
609 276
627 276
627 292
631 292
12 2 6 0 0 8320 0 10 1 0 0 5
486 313
486 348
632 348
632 310
631 310
0 5 7 0 0 8192 0 0 9 12 0 3
532 293
532 294
539 294
0 2 7 0 0 0 0 0 9 12 0 3
532 269
532 267
539 267
0 1 7 0 0 0 0 0 9 12 0 3
532 259
532 258
539 258
0 6 7 0 0 4224 0 0 9 16 0 4
405 238
532 238
532 303
539 303
0 1 7 0 0 0 0 0 10 16 0 3
407 261
407 259
416 259
0 2 7 0 0 0 0 0 10 16 0 3
407 269
407 268
416 268
0 5 7 0 0 0 0 0 10 16 0 3
407 294
407 295
416 295
1 6 7 0 0 0 0 3 10 0 0 4
375 238
407 238
407 304
416 304
0 1 8 0 0 8192 0 0 4 23 0 5
493 268
513 268
513 197
575 197
575 173
0 1 9 0 0 4224 0 0 5 22 0 4
521 276
521 203
551 203
551 174
0 1 10 0 0 4096 0 0 6 21 0 2
527 226
527 175
11 1 11 0 0 12416 0 9 7 0 0 5
603 303
621 303
621 212
502 212
502 175
9 7 10 0 0 16512 0 9 9 0 0 6
603 267
613 267
613 223
527 223
527 312
533 312
11 3 9 0 0 0 0 10 9 0 0 4
480 304
521 304
521 276
533 276
9 7 8 0 0 12416 0 10 10 0 0 6
480 268
494 268
494 222
401 222
401 313
410 313
3 3 12 0 0 4224 0 8 10 0 0 2
335 277
410 277
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
