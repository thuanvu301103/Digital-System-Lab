CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
300 130 15 200 10
336 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
336 80 1534 795
9437202 0
0
6 Title:
5 Name:
0
0
0
6
14 Logic Display~
6 431 213 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8193 0 0
2
44767.7 0
0
14 Logic Display~
6 408 213 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3917 0 0
2
44767.7 0
0
2 +V
167 238 297 0 1 3
0 4
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5723 0 0
2
44767.7 0
0
10 2-In XNOR~
219 419 293 0 3 22
0 2 3 5
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
5590 0 0
2
44767.7 0
0
7 Pulser~
4 194 247 0 10 12
0 8 9 10 7 0 0 10 10 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8500 0 0
2
44767.6 0
0
6 74LS74
17 335 264 0 12 25
0 7 6 4 4 7 5 4 4 3
6 2 11
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 0 0 0 0
1 U
4832 0 0
2
44767.6 0
0
12
0 1 2 0 0 4224 0 0 2 8 0 3
390 284
390 231
408 231
0 1 3 0 0 4096 0 0 1 9 0 3
382 237
431 237
431 231
4 0 4 0 0 4096 0 6 0 0 6 2
297 255
264 255
7 0 4 0 0 0 0 6 0 0 6 2
297 291
264 291
8 0 4 0 0 0 0 6 0 0 6 2
297 300
264 300
3 1 4 0 0 8320 0 6 3 0 0 4
297 246
264 246
264 306
238 306
3 6 5 0 0 8320 0 4 6 0 0 5
458 293
458 327
286 327
286 282
303 282
11 1 2 0 0 0 0 6 4 0 0 3
367 282
367 284
403 284
9 2 3 0 0 8320 0 6 4 0 0 4
367 237
382 237
382 302
403 302
10 2 6 0 0 8320 0 6 6 0 0 4
373 246
373 198
303 198
303 237
0 5 7 0 0 8320 0 0 6 12 0 3
250 247
250 273
303 273
4 1 7 0 0 0 0 5 6 0 0 4
224 247
250 247
250 228
303 228
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
