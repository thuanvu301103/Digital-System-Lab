CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 60 6 200 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
176 438 1534 795
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 303 217 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3104 0 0
2
44767.9 0
0
13 Logic Switch~
5 269 220 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5413 0 0
2
44767.9 0
0
13 Logic Switch~
5 237 220 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3503 0 0
2
44767.9 0
0
13 Logic Switch~
5 239 316 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3646 0 0
2
44767.9 0
0
13 Logic Switch~
5 271 316 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3631 0 0
2
44767.9 0
0
13 Logic Switch~
5 302 316 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
638 0 0
2
44767.9 0
0
14 Logic Display~
6 429 220 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6641 0 0
2
44767.9 0
0
14 Logic Display~
6 450 220 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
896 0 0
2
44767.9 0
0
14 Logic Display~
6 471 220 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6895 0 0
2
44767.9 0
0
14 Logic Display~
6 492 219 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8482 0 0
2
44767.9 0
0
14 Logic Display~
6 513 219 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
790 0 0
2
44767.9 0
0
14 Logic Display~
6 534 219 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
338 0 0
2
44767.9 0
0
14 Logic Display~
6 554 219 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
439 0 0
2
44767.9 0
0
14 Logic Display~
6 575 218 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
730 0 0
2
44767.9 0
0
7 74LS138
19 368 250 0 14 29
0 2 3 4 5 6 7 15 14 8
9 10 11 12 13
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
3377 0 0
2
44767.9 0
0
14
1 1 2 0 0 8320 0 3 15 0 0 5
249 220
249 249
328 249
328 223
336 223
1 2 3 0 0 8320 0 2 15 0 0 3
281 220
281 232
336 232
1 3 4 0 0 4224 0 1 15 0 0 3
315 217
315 241
336 241
1 4 5 0 0 8320 0 4 15 0 0 3
251 316
251 268
336 268
1 5 6 0 0 8320 0 5 15 0 0 3
283 316
283 277
330 277
1 6 7 0 0 8320 0 6 15 0 0 3
314 316
330 316
330 286
9 1 8 0 0 12416 0 15 9 0 0 5
406 241
412 241
412 246
471 246
471 238
10 1 9 0 0 4224 0 15 10 0 0 3
406 250
492 250
492 237
11 1 10 0 0 4224 0 15 11 0 0 3
406 259
513 259
513 237
12 1 11 0 0 4224 0 15 12 0 0 3
406 268
534 268
534 237
13 1 12 0 0 4224 0 15 13 0 0 3
406 277
554 277
554 237
14 1 13 0 0 4224 0 15 14 0 0 3
406 286
575 286
575 236
8 1 14 0 0 12416 0 15 8 0 0 5
406 232
416 232
416 243
450 243
450 238
7 1 15 0 0 8320 0 15 7 0 0 4
406 223
420 223
420 238
429 238
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
