CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 6 200 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
176 438 1534 795
9437202 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 293 287 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3626 0 0
2
44768 0
0
13 Logic Switch~
5 264 287 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
890 0 0
2
44768 0
0
13 Logic Switch~
5 232 286 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8835 0 0
2
44768 0
0
13 Logic Switch~
5 199 286 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9393 0 0
2
44768 0
0
13 Logic Switch~
5 167 288 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
335 0 0
2
44768 0
0
13 Logic Switch~
5 137 289 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9133 0 0
2
44768 0
0
13 Logic Switch~
5 108 290 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
792 0 0
2
44768 0
0
13 Logic Switch~
5 78 290 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
98 0 0
2
44768 0
0
13 Logic Switch~
5 293 199 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8789 0 0
2
44768 0
0
13 Logic Switch~
5 261 200 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3569 0 0
2
44768 0
0
13 Logic Switch~
5 231 200 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5300 0 0
2
44768 0
0
13 Logic Switch~
5 200 200 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3232 0 0
2
44768 0
0
13 Logic Switch~
5 171 201 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
349 0 0
2
44768 0
0
13 Logic Switch~
5 141 201 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4364 0 0
2
44768 0
0
13 Logic Switch~
5 111 202 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
936 0 0
2
44768 0
0
13 Logic Switch~
5 79 202 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6514 0 0
2
44768 0
0
14 Logic Display~
6 564 366 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3508 0 0
2
44768 0
0
14 Logic Display~
6 564 333 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3884 0 0
2
44768 0
0
14 Logic Display~
6 564 299 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9638 0 0
2
44768 0
0
7 Ground~
168 448 126 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5692 0 0
2
44768 0
0
2 +V
167 398 156 0 1 3
0 22
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3488 0 0
2
44768 0
0
6 74LS85
106 481 316 0 14 29
0 5 6 7 8 13 14 3 15 25
24 23 21 20 19
0
0 0 5104 0
5 74F85
-18 -52 17 -44
2 U2
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
3908 0 0
2
44768 0
0
6 74LS85
106 354 273 0 14 29
0 9 10 11 12 4 16 17 18 2
22 2 25 24 23
0
0 0 5104 0
5 74F85
-18 -52 17 -44
2 U1
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
6551 0 0
2
44768 0
0
26
1 7 3 0 0 8320 0 6 22 0 0 3
149 289
149 343
449 343
1 5 4 0 0 8320 0 4 23 0 0 5
211 286
211 320
314 320
314 282
322 282
1 1 5 0 0 8320 0 16 22 0 0 4
91 202
91 160
449 160
449 289
1 2 6 0 0 8320 0 15 22 0 0 5
123 202
123 168
443 168
443 298
449 298
1 3 7 0 0 8320 0 14 22 0 0 5
153 201
153 172
438 172
438 307
449 307
1 4 8 0 0 8320 0 13 22 0 0 5
183 201
183 164
434 164
434 316
449 316
1 1 9 0 0 8320 0 12 23 0 0 3
212 200
212 246
322 246
1 2 10 0 0 8320 0 11 23 0 0 3
243 200
243 255
322 255
1 3 11 0 0 12416 0 10 23 0 0 5
273 200
273 210
310 210
310 264
322 264
1 4 12 0 0 4224 0 9 23 0 0 3
305 199
305 273
322 273
1 5 13 0 0 8320 0 8 22 0 0 3
90 290
90 325
449 325
1 6 14 0 0 8320 0 7 22 0 0 3
120 290
120 334
449 334
1 0 3 0 0 128 0 6 0 0 0 3
149 289
149 292
147 292
1 8 15 0 0 8320 0 5 22 0 0 3
179 288
179 352
449 352
1 6 16 0 0 8320 0 3 23 0 0 4
244 286
244 315
322 315
322 291
1 7 17 0 0 8320 0 2 23 0 0 3
276 287
276 300
322 300
1 8 18 0 0 4224 0 1 23 0 0 3
305 287
305 309
322 309
14 1 19 0 0 8320 0 22 17 0 0 3
513 352
513 384
564 384
1 13 20 0 0 4224 0 18 22 0 0 4
564 351
533 351
533 343
513 343
1 12 21 0 0 4224 0 19 22 0 0 3
564 317
513 317
513 334
9 0 2 0 0 4096 0 23 0 0 22 2
386 246
405 246
1 11 2 0 0 8320 0 20 23 0 0 4
448 120
405 120
405 264
386 264
10 1 22 0 0 8320 0 23 21 0 0 3
386 255
398 255
398 165
14 11 23 0 0 12416 0 23 22 0 0 6
386 309
428 309
428 236
540 236
540 307
513 307
13 10 24 0 0 12416 0 23 22 0 0 6
386 300
423 300
423 244
533 244
533 298
513 298
12 9 25 0 0 12416 0 23 22 0 0 6
386 291
413 291
413 250
526 250
526 289
513 289
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
