CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
160 180 30 380 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 176 272 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8665 0 0
2
44767.7 3
0
13 Logic Switch~
5 210 272 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6236 0 0
2
44767.7 2
0
13 Logic Switch~
5 243 272 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6919 0 0
2
44767.7 1
0
13 Logic Switch~
5 279 272 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9681 0 0
2
44767.7 0
0
13 Logic Switch~
5 279 239 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3121 0 0
2
44767.7 0
0
13 Logic Switch~
5 244 238 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4121 0 0
2
44767.7 0
0
13 Logic Switch~
5 211 238 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3350 0 0
2
44767.7 0
0
13 Logic Switch~
5 177 238 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7475 0 0
2
44767.7 0
0
13 Logic Switch~
5 302 331 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 CIN
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4379 0 0
2
44767.7 0
0
14 Logic Display~
6 422 320 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4311 0 0
2
44767.7 0
0
14 Logic Display~
6 496 267 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6388 0 0
2
44767.7 0
0
14 Logic Display~
6 475 267 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
327 0 0
2
44767.7 0
0
14 Logic Display~
6 453 267 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3385 0 0
2
44767.7 0
0
14 Logic Display~
6 431 267 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6355 0 0
2
44767.7 0
0
6 74LS83
105 362 282 0 14 29
0 9 8 7 6 5 4 3 2 10
15 14 13 12 11
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3852 0 0
2
44767.7 0
0
14
1 8 2 0 0 8320 0 4 15 0 0 3
291 272
291 309
330 309
1 7 3 0 0 8320 0 3 15 0 0 3
255 272
255 300
330 300
1 6 4 0 0 8320 0 2 15 0 0 3
222 272
222 291
330 291
1 5 5 0 0 8320 0 1 15 0 0 3
188 272
188 282
330 282
1 4 6 0 0 12416 0 5 15 0 0 5
291 239
291 189
317 189
317 273
330 273
1 3 7 0 0 12416 0 6 15 0 0 5
256 238
256 194
322 194
322 264
330 264
1 2 8 0 0 8320 0 7 15 0 0 5
223 238
223 200
326 200
326 255
330 255
1 1 9 0 0 8320 0 8 15 0 0 4
189 238
189 208
330 208
330 246
1 9 10 0 0 4224 0 9 15 0 0 3
314 331
330 331
330 327
14 1 11 0 0 12416 0 15 10 0 0 4
394 327
402 327
402 338
422 338
13 1 12 0 0 12416 0 15 11 0 0 5
394 300
404 300
404 303
496 303
496 285
12 1 13 0 0 12416 0 15 12 0 0 5
394 291
408 291
408 297
475 297
475 285
11 1 14 0 0 12416 0 15 13 0 0 5
394 282
412 282
412 289
453 289
453 285
10 1 15 0 0 4224 0 15 14 0 0 4
394 273
417 273
417 285
431 285
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
