CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 100 6 270 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
176 438 1534 795
9437202 0
0
6 Title:
5 Name:
0
0
0
12
5 4081~
219 780 238 0 3 22
0 3 2 6
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
5751 0 0
2
44767.9 0
0
5 4071~
219 723 277 0 3 22
0 5 4 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3301 0 0
2
44767.9 0
0
14 Logic Display~
6 710 125 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 D
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7261 0 0
2
44767.9 0
0
14 Logic Display~
6 621 125 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9606 0 0
2
44767.9 0
0
14 Logic Display~
6 547 127 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3754 0 0
2
44767.8 0
0
14 Logic Display~
6 470 128 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9985 0 0
2
44767.8 0
0
2 +V
167 388 168 0 1 3
0 11
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5936 0 0
2
44767.8 0
0
5 4027~
219 664 261 0 7 32
0 13 14 7 15 6 16 3
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3234 0 0
2
44767.8 0
0
5 4027~
219 589 261 0 7 32
0 17 18 8 19 6 7 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
5571 0 0
2
44767.8 0
0
5 4027~
219 517 261 0 7 32
0 20 21 9 22 6 8 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7116 0 0
2
44767.8 0
0
5 4027~
219 440 260 0 7 32
0 23 11 12 11 6 9 10
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
62 0 0
2
44767.8 0
0
7 Pulser~
4 356 241 0 10 12
0 24 25 12 26 0 0 10 10 10
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3402 0 0
2
44767.7 0
0
18
3 2 2 0 0 4224 0 2 1 0 0 2
756 277
756 247
0 1 3 0 0 4224 0 0 1 9 0 3
710 183
756 183
756 229
0 2 4 0 0 8320 0 0 2 14 0 3
547 225
547 286
710 286
0 1 5 0 0 8320 0 0 2 10 0 3
621 225
621 268
710 268
0 5 6 0 0 8192 0 0 8 8 0 3
663 309
664 309
664 267
0 5 6 0 0 0 0 0 9 8 0 3
590 309
589 309
589 267
0 5 6 0 0 0 0 0 10 8 0 3
516 309
517 309
517 267
3 5 6 0 0 8320 0 1 11 0 0 4
801 238
801 309
440 309
440 266
1 7 3 0 0 4224 0 3 8 0 0 3
710 143
710 225
688 225
1 7 5 0 0 128 0 4 9 0 0 3
621 143
621 225
613 225
6 3 7 0 0 12416 0 9 8 0 0 4
619 243
629 243
629 234
640 234
6 3 8 0 0 4224 0 10 9 0 0 4
547 243
557 243
557 234
565 234
6 3 9 0 0 12416 0 11 10 0 0 4
470 242
480 242
480 234
493 234
1 7 4 0 0 128 0 5 10 0 0 3
547 145
547 225
541 225
1 7 10 0 0 4224 0 6 11 0 0 3
470 146
470 224
464 224
0 2 11 0 0 8192 0 0 11 17 0 3
408 223
408 224
416 224
1 4 11 0 0 12416 0 7 11 0 0 5
388 177
388 196
408 196
408 242
416 242
3 3 12 0 0 8320 0 12 11 0 0 3
380 232
380 233
416 233
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
