CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 150 15 310 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 60 310 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5949 0 0
2
44767.7 0
0
13 Logic Switch~
5 60 264 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
31 0 0
2
44767.7 0
0
13 Logic Switch~
5 59 226 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3515 0 0
2
44767.7 0
0
14 Logic Display~
6 460 278 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4916 0 0
2
44767.7 0
0
14 Logic Display~
6 404 210 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9329 0 0
2
44767.7 0
0
5 4071~
219 393 297 0 3 22
0 4 5 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3773 0 0
2
44767.7 0
0
5 4081~
219 302 296 0 3 22
0 7 6 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3544 0 0
2
44767.7 0
0
5 4081~
219 177 301 0 3 22
0 9 8 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
4373 0 0
2
44767.7 0
0
5 4030~
219 298 231 0 3 22
0 7 6 3
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3405 0 0
2
44767.7 0
0
5 4030~
219 173 234 0 3 22
0 9 8 7
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
327 0 0
2
44767.7 0
0
12
3 1 2 0 0 8320 0 6 4 0 0 3
426 297
426 296
460 296
3 1 3 0 0 4224 0 9 5 0 0 3
331 231
404 231
404 228
3 1 4 0 0 8320 0 7 6 0 0 3
323 296
323 288
380 288
3 2 5 0 0 12416 0 8 6 0 0 6
198 301
221 301
221 318
350 318
350 306
380 306
0 2 6 0 0 4096 0 0 7 7 0 3
259 240
259 305
278 305
0 1 7 0 0 4224 0 0 7 8 0 3
272 222
272 287
278 287
1 2 6 0 0 12416 0 1 9 0 0 6
72 310
109 310
109 332
249 332
249 240
282 240
3 1 7 0 0 0 0 10 9 0 0 4
206 234
236 234
236 222
282 222
0 2 8 0 0 4224 0 0 8 11 0 3
123 243
123 310
153 310
0 1 9 0 0 4096 0 0 8 12 0 3
140 225
140 292
153 292
1 2 8 0 0 0 0 2 10 0 0 4
72 264
112 264
112 243
157 243
1 1 9 0 0 8320 0 3 10 0 0 3
71 226
71 225
157 225
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
