CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 140 15 480 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
6
2 +V
167 338 267 0 1 3
0 4
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
428 0 0
2
5.9004e-315 0
0
10 2-In XNOR~
219 500 232 0 3 22
0 3 2 5
0
0 0 608 0
4 4077
-7 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
6112 0 0
2
5.9004e-315 0
0
14 Logic Display~
6 525 170 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
492 0 0
2
5.9004e-315 0
0
14 Logic Display~
6 497 170 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7418 0 0
2
5.9004e-315 0
0
7 Pulser~
4 308 209 0 10 12
0 8 9 10 7 0 0 10 10 1
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7724 0 0
2
5.9004e-315 0
0
6 74LS74
17 422 230 0 12 25
0 7 6 4 4 7 5 4 4 3
6 2 11
0
0 0 4832 0
6 74LS74
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 1 0 0 0
1 U
4426 0 0
2
5.9004e-315 0
0
12
0 1 2 0 0 4224 0 0 4 8 0 3
479 241
479 188
497 188
0 1 3 0 0 4224 0 0 3 9 0 3
470 203
525 203
525 188
8 0 4 0 0 4096 0 6 0 0 6 2
384 266
367 266
7 0 4 0 0 0 0 6 0 0 6 2
384 257
367 257
4 0 4 0 0 0 0 6 0 0 6 2
384 221
367 221
3 1 4 0 0 8320 0 6 1 0 0 4
384 212
367 212
367 276
338 276
3 6 5 0 0 8320 0 2 6 0 0 5
539 232
539 282
380 282
380 248
390 248
11 2 2 0 0 0 0 6 2 0 0 4
454 248
470 248
470 241
484 241
9 1 3 0 0 0 0 6 2 0 0 4
454 203
470 203
470 223
484 223
10 2 6 0 0 8320 0 6 6 0 0 5
460 212
460 165
381 165
381 203
390 203
0 4 7 0 0 4096 0 0 5 12 0 2
352 209
338 209
1 5 7 0 0 8320 0 6 6 0 0 4
390 194
352 194
352 239
390 239
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
